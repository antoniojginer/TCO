* C:\Users\Antonio Jose\Documents\UPV\TCO\practicas\pract4.sch

* Schematics Version 9.1 - Web Update 1
* Tue May 29 20:49:58 2018



** Analysis setup **
.tran 1n 1u
.LIB "C:\Users\Antonio Jose\Documents\UPV\TCO\practicas\pract4.lib"
.STMLIB "pract4.stl"


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "pract4.net"
.INC "pract4.als"


.probe


.END
