* C:\Users\Antonio Jose\Documents\UPV\TCO\practicas\Schematic1.sch

* Schematics Version 9.1 - Web Update 1
* Tue May 29 22:33:52 2018



** Analysis setup **
.DC LIN V_V1 0 5 0.01 
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "Schematic1.net"
.INC "Schematic1.als"


.probe


.END
